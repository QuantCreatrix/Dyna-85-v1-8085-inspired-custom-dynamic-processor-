// controlStates.vh - Control Unit State Definitions

// Main states
`define STATE_FETCH     4'b0000
`define STATE_DECODE    4'b0001

// Single-byte instruction states
`define STATE_MOV_EXEC  4'b0010
