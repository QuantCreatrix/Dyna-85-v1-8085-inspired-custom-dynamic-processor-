// registers.vh - Register Definitions

// General Purpose Registers
`define REG_A       3'b000
`define REG_B       3'b001
`define REG_C       3'b010
`define REG_D       3'b011
`define REG_E       3'b100
`define REG_H       3'b101
`define REG_L       3'b110